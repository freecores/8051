
///
/// created by p8051Rom.exe
/// author: Simon Teran (simont@opencores.org)
///
/// source file: D:\verilog\oc8051\test\TMP\Negcnt.ihx
/// date: 6.6.02
/// time: 22:02:17
///

module oc8051_rom (rst, clk, addr, ea_int, data1, data2, data3);

parameter INT_ROM_WID= 15;

input rst, clk;
input [15:0] addr;
output ea_int;
output [7:0] data1, data2, data3;

reg ea_int;
reg [7:0] data1, data2, data3;
reg [7:0] buff [65535:0];
integer i;

wire ea;

assign ea = | addr[15:INT_ROM_WID];
//assign ea_int = ! ea;

initial
begin
  for (i=0; i<65536; i=i+1)
    buff [i] = 8'h00;
  $readmemh("../src/oc8051_rom.in", buff);
end

always @(posedge clk or posedge rst)
 if (rst)
   ea_int <= #1 1'b1;
  else ea_int <= #1 !ea;

always @(posedge clk)
begin
  data1 <= #1 buff [addr];
  data2 <= #1 buff [addr+1];
  data3 <= #1 buff [addr+2];
end

endmodule


